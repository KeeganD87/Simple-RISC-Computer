module rotate_left(
	output [31:0] R,
	input [31:0] A, B
);
	wire [4:0] N;
	assign N = A % 32;
	assign R =  (N == 31)?{B[0:0], B[31:1]}:
				   (N == 30)?{B[1:0], B[31:2]}:
				   (N == 29)?{B[2:0], B[31:3]}:
					(N == 28)?{B[3:0], B[31:4]}:
					(N == 27)?{B[4:0], B[31:5]}:
					(N == 26)?{B[5:0], B[31:6]}:
					(N == 25)?{B[6:0], B[31:7]}:
					(N == 24)?{B[7:0], B[31:8]}:
					(N == 23)?{B[8:0], B[31:9]}:
					(N == 22)?{B[9:0], B[31:10]}:
					(N == 21)?{B[10:0], B[31:11]}:
					(N == 20)?{B[11:0], B[31:12]}:
					(N == 19)?{B[12:0], B[31:13]}:
					(N == 18)?{B[13:0], B[31:14]}:
					(N == 17)?{B[14:0], B[31:15]}:
					(N == 16)?{B[15:0], B[31:16]}:
					(N == 15)?{B[16:0], B[31:17]}:
					(N == 14)?{B[17:0], B[31:18]}:
					(N == 13)?{B[18:0], B[31:19]}:
					(N == 12)?{B[19:0], B[31:20]}:
					(N == 11)?{B[20:0], B[31:21]}:
					(N == 10)?{B[21:0], B[31:22]}:
					(N == 9)?{B[22:0], B[31:23]}:
					(N == 8)?{B[23:0], B[31:24]}:
					(N == 7)?{B[24:0], B[31:25]}:
					(N == 6)?{B[25:0], B[31:26]}:
					(N == 5)?{B[26:0], B[31:27]}:
					(N == 4)?{B[27:0], B[31:28]}:
					(N == 3)?{B[28:0], B[31:29]}:
					(N == 2)?{B[29:0], B[31:30]}:
					(N == 1)?{B[30:0], B[31:31]}:
					B[31:0];

endmodule

 module rotate_right(
	output [31:0] R,
	input [31:0] A, B
 );
	wire [4:0] N;
	assign N = A % 32;
	assign R =  (N == 31)?{B[30:0], B[31:31]}:
					(N == 30)?{B[29:0], B[31:30]}:
					(N == 29)?{B[28:0], B[31:29]}:
					(N == 28)?{B[27:0], B[31:28]}:
					(N == 27)?{B[26:0], B[31:27]}:
					(N == 26)?{B[25:0], B[31:26]}:
					(N == 25)?{B[24:0], B[31:25]}:
					(N == 24)?{B[23:0], B[31:24]}:
					(N == 23)?{B[22:0], B[31:23]}:
					(N == 22)?{B[21:0], B[31:22]}:
					(N == 21)?{B[20:0], B[31:21]}:
					(N == 20)?{B[19:0], B[31:20]}:
					(N == 19)?{B[18:0], B[31:19]}:
					(N == 18)?{B[17:0], B[31:18]}:
					(N == 17)?{B[16:0], B[31:17]}:
					(N == 16)?{B[15:0], B[31:16]}:
					(N == 15)?{B[14:0], B[31:15]}:
					(N == 14)?{B[13:0], B[31:14]}:
					(N == 13)?{B[12:0], B[31:13]}:
					(N == 12)?{B[11:0], B[31:12]}:
					(N == 11)?{B[10:0], B[31:11]}:
					(N == 10)?{B[9:0], B[31:10]}:
					(N == 9)?{B[8:0], B[31:9]}:
					(N == 8)?{B[7:0], B[31:8]}:
					(N == 7)?{B[6:0], B[31:7]}:
					(N == 6)?{B[5:0], B[31:6]}:
					(N == 5)?{B[4:0], B[31:5]}:
					(N == 4)?{B[3:0], B[31:4]}:
					(N == 3)?{B[2:0], B[31:3]}:
					(N == 2)?{B[1:0], B[31:2]}:
					(N == 1)?{B[0:0], B[31:1]}:
					B[31:0];
					
endmodule
